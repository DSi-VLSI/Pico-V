////////////////////////////////////////////////////////////////////////////////////////////////////
// 
//  File:        tb_template.sv
//  Author:      <Your Name>
//  Created:     <Date>
//  Description: A general-purpose SystemVerilog testbench template. This template provides a
//               structured starting point for verifying a Design Under Test (DUT).
// 
////////////////////////////////////////////////////////////////////////////////////////////////////

module tb_template;

  initial begin
    $display("Hello World!");
    $finish;
  end

endmodule